
interface pe_intf;
	// All signals declaration which present inside the DUT
	bit a0;
	bit a1;
	bit a2;
	bit a3;
	bit y0;
	bit y1;
	bit v;
	
	// Declaration of clocking bloks 
	// Declaration of the modports
endinterface